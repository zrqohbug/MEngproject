`timescale 1ns / 1ps
module tb
#(
	parameter data_size = 8
);


 // Inputs
 reg clk;
 reg reset;
 reg [data_size-1:0] a1;
 reg [data_size-1:0] a2;
 reg [data_size-1:0] b1;
 reg [data_size-1:0] b2;


 // Outputs
 wire [2*data_size-1:0] c1;
 wire [2*data_size-1:0] c2;
 wire [2*data_size-1:0] c3;
 wire [2*data_size-1:0] c4;


 // Instantiate the Unit Under Test (UUT)
  systolictop test(
  .clk(clk), 
  .reset(reset), 
  .a1(a1), 
  .a2(a2), 
  .b1(b1), 
  .b2(b2), 
  .c1(c1), 
  .c2(c2), 
  .c3(c3), 
  .c4(c4),
  .v(0),
  .x(0),
  .y(0)
 );

 initial begin
  // Initialize Inputs
  clk = 0;
  reset = 0;
  a1 = 0;
  a2 = 0;
  b1 = 0;
  b2 = 0;


  // assume we have a matrix A
  //[1,2,3,4,5,6,7,8]
  //[2,3,4,5,6,7,8,1]
  //[3,4,5,6,7,8,1,2]
  //[4,5,6,7,8,1,2,3]
  //[5,6,7,8,1,2,3,4]
  //[6,7,8,1,2,3,4,5]
  //[7,8,1,2,3,4,5,6]
  //[8,1,2,3,4,5,6,7]

    // assume we have a matrix B
  //[0,1,2,3,4,5,6,7]
  //[1,2,3,4,5,6,7,0]
  //[2,3,4,5,6,7,0,1]
  //[3,4,5,6,7,0,1,2]
  //[4,5,6,7,0,1,2,3]
  //[5,6,7,0,1,2,3,4]
  //[6,7,0,1,2,3,4,5]
  //[7,0,1,2,3,4,5,6]


  // Wait 100 ns for global reset to finish
  #5 reset = 1;
  #5 reset = 0;

  #10; a1 = 1; a2 = 0;  b1 = 0; b2 = 0; 

  #10; a1 = 2; a2 = 2;  b1 = 1; b2 = 1;
  #10; a1 = 3; a2 = 3;  b1 = 2; b2 = 2; 
  #10; a1 = 4; a2 = 4;  b1 = 3; b2 = 3; 
  #10; a1 = 5; a2 = 5;  b1 = 4; b2 = 4; 
  #10; a1 = 6; a2 = 6;  b1 = 5; b2 = 5; 
  #10; a1 = 7; a2 = 7;  b1 = 6; b2 = 6; 
  #10; a1 = 8; a2 = 8;  b1 = 7; b2 = 7;

  #10; a1 = 1; a2 = 1;  b1 = 2; b2 = 0;

  #10; a1 = 2; a2 = 2;  b1 = 3; b2 = 3; 
  #10; a1 = 3; a2 = 3;  b1 = 4; b2 = 4;
  #10; a1 = 4; a2 = 4;  b1 = 5; b2 = 5; 
  #10; a1 = 5; a2 = 5;  b1 = 6; b2 = 6; 
  #10; a1 = 6; a2 = 6;  b1 = 7; b2 = 7; 
  #10; a1 = 7; a2 = 7;  b1 = 0; b2 = 0;
  #10; a1 = 8; a2 = 8;  b1 = 1; b2 = 1; 

  #10; a1 = 1; a2 = 1;  b1 = 4; b2 = 2;

  #10; a1 = 2; a2 = 2;  b1 = 5; b2 = 5; 
  #10; a1 = 3; a2 = 3;  b1 = 6; b2 = 6;
  #10; a1 = 4; a2 = 4;  b1 = 7; b2 = 7; 
  #10; a1 = 5; a2 = 5;  b1 = 0; b2 = 0; 
  #10; a1 = 6; a2 = 6;  b1 = 1; b2 = 1; 
  #10; a1 = 7; a2 = 7;  b1 = 2; b2 = 2;
  #10; a1 = 8; a2 = 8;  b1 = 3; b2 = 3; 

  #10; a1 = 1; a2 = 1;  b1 = 6; b2 = 4;

  #10; a1 = 2; a2 = 2;  b1 = 7; b2 = 7; 
  #10; a1 = 3; a2 = 3;  b1 = 0; b2 = 0;
  #10; a1 = 4; a2 = 4;  b1 = 1; b2 = 1; 
  #10; a1 = 5; a2 = 5;  b1 = 2; b2 = 2; 
  #10; a1 = 6; a2 = 6;  b1 = 3; b2 = 3; 
  #10; a1 = 7; a2 = 7;  b1 = 4; b2 = 4;
  #10; a1 = 8; a2 = 8;  b1 = 5; b2 = 5; 

  #10; a1 = 3; a2 = 1;  b1 = 0; b2 = 6;

//////////////////////////////////////////
/////// A1 and A2   //////////////////////
//////////////////////////////////////////


  #10; a1 = 4; a2 = 4;  b1 = 1; b2 = 1;
  #10; a1 = 5; a2 = 5;  b1 = 2; b2 = 2; 
  #10; a1 = 6; a2 = 6;  b1 = 3; b2 = 3; 
  #10; a1 = 7; a2 = 7;  b1 = 4; b2 = 4; 
  #10; a1 = 8; a2 = 8;  b1 = 5; b2 = 5; 
  #10; a1 = 1; a2 = 1;  b1 = 6; b2 = 6; 
  #10; a1 = 2; a2 = 2;  b1 = 7; b2 = 7;

  #10; a1 = 3; a2 = 3;  b1 = 2; b2 = 0;

  #10; a1 = 4; a2 = 4;  b1 = 3; b2 = 3; 
  #10; a1 = 5; a2 = 5;  b1 = 4; b2 = 4;
  #10; a1 = 6; a2 = 6;  b1 = 5; b2 = 5; 
  #10; a1 = 7; a2 = 7;  b1 = 6; b2 = 6; 
  #10; a1 = 8; a2 = 8;  b1 = 7; b2 = 7; 
  #10; a1 = 1; a2 = 1;  b1 = 0; b2 = 0;
  #10; a1 = 2; a2 = 2;  b1 = 1; b2 = 1; 

  #10; a1 = 3; a2 = 3;  b1 = 4; b2 = 2;

  #10; a1 = 4; a2 = 4;  b1 = 5; b2 = 5; 
  #10; a1 = 5; a2 = 5;  b1 = 6; b2 = 6;
  #10; a1 = 6; a2 = 6;  b1 = 7; b2 = 7; 
  #10; a1 = 7; a2 = 7;  b1 = 0; b2 = 0; 
  #10; a1 = 8; a2 = 8;  b1 = 1; b2 = 1; 
  #10; a1 = 1; a2 = 1;  b1 = 2; b2 = 2;
  #10; a1 = 2; a2 = 2;  b1 = 3; b2 = 3; 

  #10; a1 = 3; a2 = 3;  b1 = 6; b2 = 4;

  #10; a1 = 4; a2 = 4;  b1 = 7; b2 = 7; 
  #10; a1 = 5; a2 = 5;  b1 = 0; b2 = 0;
  #10; a1 = 6; a2 = 6;  b1 = 1; b2 = 1; 
  #10; a1 = 7; a2 = 7;  b1 = 2; b2 = 2; 
  #10; a1 = 8; a2 = 8;  b1 = 3; b2 = 3; 
  #10; a1 = 1; a2 = 1;  b1 = 4; b2 = 4;
  #10; a1 = 2; a2 = 2;  b1 = 5; b2 = 5; 

  #10; a1 = 5; a2 = 3;  b1 = 0; b2 = 6;


//////////////////////////////////////////
/////// A3 and A4   //////////////////////
//////////////////////////////////////////


  #10; a1 = 6; a2 = 6;  b1 = 1; b2 = 1;
  #10; a1 = 7; a2 = 7;  b1 = 2; b2 = 2; 
  #10; a1 = 8; a2 = 8;  b1 = 3; b2 = 3; 
  #10; a1 = 1; a2 = 1;  b1 = 4; b2 = 4; 
  #10; a1 = 2; a2 = 2;  b1 = 5; b2 = 5; 
  #10; a1 = 3; a2 = 3;  b1 = 6; b2 = 6; 
  #10; a1 = 4; a2 = 4;  b1 = 7; b2 = 7;

  #10; a1 = 5; a2 = 5;  b1 = 2; b2 = 0;

  #10; a1 = 6; a2 = 6;  b1 = 3; b2 = 3; 
  #10; a1 = 7; a2 = 7;  b1 = 4; b2 = 4;
  #10; a1 = 8; a2 = 8;  b1 = 5; b2 = 5; 
  #10; a1 = 1; a2 = 1;  b1 = 6; b2 = 6; 
  #10; a1 = 2; a2 = 2;  b1 = 7; b2 = 7; 
  #10; a1 = 3; a2 = 3;  b1 = 0; b2 = 0;
  #10; a1 = 4; a2 = 4;  b1 = 1; b2 = 1; 

  #10; a1 = 3; a2 = 3;  b1 = 4; b2 = 2;

  #10; a1 = 4; a2 = 4;  b1 = 5; b2 = 5; 
  #10; a1 = 5; a2 = 5;  b1 = 6; b2 = 6;
  #10; a1 = 6; a2 = 6;  b1 = 7; b2 = 7; 
  #10; a1 = 7; a2 = 7;  b1 = 0; b2 = 0; 
  #10; a1 = 8; a2 = 8;  b1 = 1; b2 = 1; 
  #10; a1 = 1; a2 = 1;  b1 = 2; b2 = 2;
  #10; a1 = 2; a2 = 2;  b1 = 3; b2 = 3; 

  #10; a1 = 3; a2 = 3;  b1 = 6; b2 = 4;

  #10; a1 = 4; a2 = 4;  b1 = 7; b2 = 7; 
  #10; a1 = 5; a2 = 5;  b1 = 0; b2 = 0;
  #10; a1 = 6; a2 = 6;  b1 = 1; b2 = 1; 
  #10; a1 = 7; a2 = 7;  b1 = 2; b2 = 2; 
  #10; a1 = 8; a2 = 8;  b1 = 3; b2 = 3; 
  #10; a1 = 1; a2 = 1;  b1 = 4; b2 = 4;
  #10; a1 = 2; a2 = 2;  b1 = 5; b2 = 5; 

  #10; a1 = 3; a2 = 3;  b1 = 4; b2 = 6;

////////////////////////////////////////////////////////////////////////////
  #10; a1 = 1 ; a2 = 0;  b1 = 0; b2 = 0; 

  for (i = 0; i <= 7; i = i+2)
  	for (j = 0; j <= 7; j = j+2)
  	{
  		  #10; a1 = i + 2 ; a2 = i + 2;  b1 = (j + 1) % 8; b2 = (j + 1) % 8; 
   		  #10; a1 = i + 3 ; a2 = i + 3;  b1 = (j + 2) % 8; b2 = (j + 2) % 8; 
   		  #10; a1 = i + 4 ; a2 = i + 4;  b1 = (j + 3) % 8; b2 = (j + 3) % 8; 
   		  #10; a1 = i + 5 ; a2 = i + 5;  b1 = (j + 4) % 8; b2 = (j + 4) % 8; 
  		  #10; a1 = i + 6 ; a2 = i + 6;  b1 = (j + 5) % 8; b2 = (j + 5) % 8; 
  		  #10; a1 = i + 7 ; a2 = i + 7;  b1 = (j + 6) % 8; b2 = (j + 6) % 8; 
  		  #10; a1 = i + 8 ; a2 = i + 8;  b1 = (j + 7) % 8; b2 = (j + 7) % 8; 
  		  if (j != 6)
  		  	#10; a1 = i + 1 ; a2 = i + 1;  b1 = (j + 2) % 8; b2 = j;
  		  else if (i != 6)
  		  	#10; a1 = i + 3 ; a2 = i + 1;  b1 = (j + 2) % 8; b2 = j; 
  		  else
  		    #10; a1 = 0 ; a2 = i + 1;  b1 = (j + 2) % 8; b2 = j;  		  	 
  	}
  #100;
  $stop;

 end
 
 always begin
   #5 clk = ~clk;

 end
      
endmodule
